-------------------------------------------------------------------------------
-- coeff_rom.vhd
-- Coefficient ROM for Polyphase Channelizer
-------------------------------------------------------------------------------
-- Open Research Institute
-- Project: Polyphase Channelizer (MDT / Haifuraiya)
-- 
-- Description:
--   Stores prototype filter coefficients in fixed-point format for the 
--   polyphase filterbank. Coefficients are distributed round-robin across
--   branches (the standard polyphase decomposition):
--   
--     Original filter: h[0], h[1], h[2], h[3], h[4], h[5], h[6], h[7], ...
--     
--     Branch 0 gets: h[0], h[N], h[2N], ...  (i.e., h[0], h[4], h[8], ... for N=4)
--     Branch 1 gets: h[1], h[N+1], h[2N+1], ...  (i.e., h[1], h[5], h[9], ...)
--     Branch 2 gets: h[2], h[N+2], h[2N+2], ...
--     ...
--     Branch N-1 gets: h[N-1], h[2N-1], h[3N-1], ...
--   
--   In ROM, coefficients are stored contiguously per branch for efficient access:
--     Address 0..M-1:           Branch 0's M coefficients
--     Address M..2M-1:          Branch 1's M coefficients
--     ...
--     Address (N-1)*M..N*M-1:   Branch N-1's M coefficients
--   
--   Where N = number of channels, M = taps per branch.
--
--   The ROM is initialized from a hex file generated by the Python reference
--   implementation, allowing the same RTL to support both MDT (64 coeffs) and
--   Haifuraiya (1536 coeffs) configurations.
--
-- Target: iCE40 UltraPlus (MDT), Xilinx ZCU102 (Haifuraiya)
--
-- Resource Usage (iCE40):
--   MDT:        64 x 16-bit  = 1,024 bits  = 1 EBR (4Kb each)
--   Haifuraiya: 1536 x 16-bit = 24,576 bits = 6 EBRs
--
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity coeff_rom is
    generic (
        -- Number of channels (N)
        -- Valid: 4 (MDT), 64 (Haifuraiya)
        N_CHANNELS      : positive := 4;
        
        -- Taps per polyphase branch (M)
        -- Total taps = N_CHANNELS * TAPS_PER_BRANCH
        -- Valid: 16 (MDT: 64 total), 24 (Haifuraiya: 1536 total)
        TAPS_PER_BRANCH : positive := 16;
        
        -- Coefficient bit width (signed fixed-point)
        -- Q1.15 format: 1 sign bit, 15 fractional bits
        COEFF_WIDTH     : positive := 16;
        
        -- Address width (must equal ceil(log2(N_CHANNELS * TAPS_PER_BRANCH)))
        -- MDT: ceil(log2(64)) = 6,  Haifuraiya: ceil(log2(1536)) = 11
        ADDR_WIDTH      : positive := 6;
        
        -- Path to coefficient hex file
        -- File format: One coefficient per line, hexadecimal, MSB first
        -- Generated by: polyphase_channelizer.ipynb
        COEFF_FILE      : string := "coeffs.hex"
    );
    port (
        -- Clock
        clk     : in  std_logic;
        
        -- Address input
        -- Range: 0 to (N_CHANNELS * TAPS_PER_BRANCH - 1)
        addr    : in  std_logic_vector(ADDR_WIDTH - 1 downto 0);
        
        -- Coefficient output (signed, 1 cycle latency)
        coeff   : out std_logic_vector(COEFF_WIDTH - 1 downto 0)
    );
end entity coeff_rom;

architecture rtl of coeff_rom is

    ---------------------------------------------------------------------------
    -- Constants
    ---------------------------------------------------------------------------
    constant ROM_DEPTH : positive := N_CHANNELS * TAPS_PER_BRANCH;
    
    ---------------------------------------------------------------------------
    -- Types
    ---------------------------------------------------------------------------
    type rom_type is array (0 to ROM_DEPTH - 1) of 
        std_logic_vector(COEFF_WIDTH - 1 downto 0);
    
    -- Initialize ROM from hex file
    -- File format: One hex value per line (e.g., "7FFF" for +0.99997)
    impure function init_rom_from_file(filename : string) return rom_type is
        file rom_file     : text;
        variable rom_line : line;
        variable rom_data : rom_type;
        variable hex_val  : std_logic_vector(COEFF_WIDTH - 1 downto 0);
        variable good     : boolean;
    begin
        -- Initialize to zero in case file is short
        for i in rom_type'range loop
            rom_data(i) := (others => '0');
        end loop;
        
        -- Read coefficients from file
        file_open(rom_file, filename, read_mode);
        for i in 0 to ROM_DEPTH - 1 loop
            exit when endfile(rom_file);
            readline(rom_file, rom_line);
            hread(rom_line, hex_val, good);
            if good then
                rom_data(i) := hex_val;
            end if;
        end loop;
        file_close(rom_file);
        
        return rom_data;
    end function init_rom_from_file;
    
    ---------------------------------------------------------------------------
    -- Signals
    ---------------------------------------------------------------------------
    signal rom : rom_type := init_rom_from_file(COEFF_FILE);
    
    -- Register for output (creates single-cycle latency, helps timing)
    signal coeff_reg : std_logic_vector(COEFF_WIDTH - 1 downto 0);

begin

    ---------------------------------------------------------------------------
    -- ROM Read Process
    ---------------------------------------------------------------------------
    -- Synchronous read with registered output
    -- This coding style infers Block RAM on both iCE40 and Xilinx
    ---------------------------------------------------------------------------
    process(clk)
    begin
        if rising_edge(clk) then
            coeff_reg <= rom(to_integer(unsigned(addr)));
        end if;
    end process;
    
    -- Output assignment
    coeff <= coeff_reg;

end architecture rtl;
